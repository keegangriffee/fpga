module cl_dma_pcis_slv
(
	input clk,
	input rst_n,
	axi_bus_t.master dma_pcis_bus,
	axi_bus_t.master mem_reader_axi,
	axi_bus_t.slave ddr_a_out,
	axi_bus_t.slave ddr_b_out,
	axi_bus_t.slave ddr_c_out,
	axi_bus_t.slave ddr_d_out
);

axi_bus_t dma_pcis_bus_q();
axi_bus_t mem_reader_axi_q();

axi_bus_t ddr_a_pre();
axi_bus_t ddr_b_pre();
axi_bus_t ddr_c_pre();
axi_bus_t ddr_d_pre();

axi_bus_t ddr_a_src();
axi_bus_t ddr_b_src();
axi_bus_t ddr_d_src();

axi_bus_t ddr_a_dest();
axi_bus_t ddr_b_dest();
axi_bus_t ddr_d_dest();

// reset sync
(* dont_touch *) logic slr_sync_aresetn;
lib_pipe #(.WIDTH(1), .STAGES(4)) SLR_PIPE_RST_N (
	.clk(clk), .rst_n(1'b1),
	.in_bus(rst_n),
	.out_bus(slr_sync_aresetn)
);

axi_register_slice DMA_PCIS_BUS_REG_SLICE
(
	.aclk(clk),
	.aresetn(slr_sync_aresetn),

	.s_axi_awid    (dma_pcis_bus.awid),
	.s_axi_awaddr  (dma_pcis_bus.awaddr),
	.s_axi_awlen   (dma_pcis_bus.awlen),                                            
	.s_axi_awvalid (dma_pcis_bus.awvalid),
	.s_axi_awsize  (dma_pcis_bus.awsize),
	.s_axi_awready (dma_pcis_bus.awready),
	.s_axi_wdata   (dma_pcis_bus.wdata),
	.s_axi_wstrb   (dma_pcis_bus.wstrb),
	.s_axi_wlast   (dma_pcis_bus.wlast),
	.s_axi_wvalid  (dma_pcis_bus.wvalid),
	.s_axi_wready  (dma_pcis_bus.wready),
	.s_axi_bid     (dma_pcis_bus.bid),
	.s_axi_bresp   (dma_pcis_bus.bresp),
	.s_axi_bvalid  (dma_pcis_bus.bvalid),
	.s_axi_bready  (dma_pcis_bus.bready),
	.s_axi_arid    (dma_pcis_bus.arid),
	.s_axi_araddr  (dma_pcis_bus.araddr),
	.s_axi_arlen   (dma_pcis_bus.arlen), 
	.s_axi_arvalid (dma_pcis_bus.arvalid),
	.s_axi_arsize  (dma_pcis_bus.arsize),
	.s_axi_arready (dma_pcis_bus.arready),
	.s_axi_rid     (dma_pcis_bus.rid),
	.s_axi_rdata   (dma_pcis_bus.rdata),
	.s_axi_rresp   (dma_pcis_bus.rresp),
	.s_axi_rlast   (dma_pcis_bus.rlast),
	.s_axi_rvalid  (dma_pcis_bus.rvalid),
	.s_axi_rready  (dma_pcis_bus.rready),

	.m_axi_awid    (dma_pcis_bus_q.awid),
	.m_axi_awaddr  (dma_pcis_bus_q.awaddr), 
	.m_axi_awlen   (dma_pcis_bus_q.awlen),
	.m_axi_awvalid (dma_pcis_bus_q.awvalid),
	.m_axi_awsize  (dma_pcis_bus_q.awsize),
	.m_axi_awready (dma_pcis_bus_q.awready),
	.m_axi_wdata   (dma_pcis_bus_q.wdata),  
	.m_axi_wstrb   (dma_pcis_bus_q.wstrb),
	.m_axi_wvalid  (dma_pcis_bus_q.wvalid), 
	.m_axi_wlast   (dma_pcis_bus_q.wlast),
	.m_axi_wready  (dma_pcis_bus_q.wready), 
	.m_axi_bresp   (dma_pcis_bus_q.bresp),  
	.m_axi_bvalid  (dma_pcis_bus_q.bvalid), 
	.m_axi_bid     (dma_pcis_bus_q.bid),
	.m_axi_bready  (dma_pcis_bus_q.bready), 
	.m_axi_arid    (dma_pcis_bus_q.arid), 
	.m_axi_araddr  (dma_pcis_bus_q.araddr), 
	.m_axi_arlen   (dma_pcis_bus_q.arlen), 
	.m_axi_arsize  (dma_pcis_bus_q.arsize), 
	.m_axi_arvalid (dma_pcis_bus_q.arvalid),
	.m_axi_arready (dma_pcis_bus_q.arready),
	.m_axi_rid     (dma_pcis_bus_q.rid),  
	.m_axi_rdata   (dma_pcis_bus_q.rdata),  
	.m_axi_rresp   (dma_pcis_bus_q.rresp),  
	.m_axi_rlast   (dma_pcis_bus_q.rlast),  
	.m_axi_rvalid  (dma_pcis_bus_q.rvalid), 
	.m_axi_rready  (dma_pcis_bus_q.rready)
);

// mem reader bus reg slice
axi_register_slice MEM_READER_AXI_REG_SLICE
(
	.aclk(clk),
	.aresetn(slr_sync_aresetn),

	.s_axi_awid    (mem_reader_axi.awid),
	.s_axi_awaddr  (mem_reader_axi.awaddr),
	.s_axi_awlen   (mem_reader_axi.awlen),                                            
	.s_axi_awvalid (mem_reader_axi.awvalid),
	.s_axi_awsize  (mem_reader_axi.awsize),
	.s_axi_awready (mem_reader_axi.awready),
	.s_axi_wdata   (mem_reader_axi.wdata),
	.s_axi_wstrb   (mem_reader_axi.wstrb),
	.s_axi_wlast   (mem_reader_axi.wlast),
	.s_axi_wvalid  (mem_reader_axi.wvalid),
	.s_axi_wready  (mem_reader_axi.wready),
	.s_axi_bid     (mem_reader_axi.bid),
	.s_axi_bresp   (mem_reader_axi.bresp),
	.s_axi_bvalid  (mem_reader_axi.bvalid),
	.s_axi_bready  (mem_reader_axi.bready),
	.s_axi_arid    (mem_reader_axi.arid),
	.s_axi_araddr  (mem_reader_axi.araddr),
	.s_axi_arlen   (mem_reader_axi.arlen), 
	.s_axi_arvalid (mem_reader_axi.arvalid),
	.s_axi_arsize  (mem_reader_axi.arsize),
	.s_axi_arready (mem_reader_axi.arready),
	.s_axi_rid     (mem_reader_axi.rid),
	.s_axi_rdata   (mem_reader_axi.rdata),
	.s_axi_rresp   (mem_reader_axi.rresp),
	.s_axi_rlast   (mem_reader_axi.rlast),
	.s_axi_rvalid  (mem_reader_axi.rvalid),
	.s_axi_rready  (mem_reader_axi.rready),

	.m_axi_awid    (mem_reader_axi_q.awid),
	.m_axi_awaddr  (mem_reader_axi_q.awaddr), 
	.m_axi_awlen   (mem_reader_axi_q.awlen),
	.m_axi_awvalid (mem_reader_axi_q.awvalid),
	.m_axi_awsize  (mem_reader_axi_q.awsize),
	.m_axi_awready (mem_reader_axi_q.awready),
	.m_axi_wdata   (mem_reader_axi_q.wdata),  
	.m_axi_wstrb   (mem_reader_axi_q.wstrb),
	.m_axi_wvalid  (mem_reader_axi_q.wvalid), 
	.m_axi_wlast   (mem_reader_axi_q.wlast),
	.m_axi_wready  (mem_reader_axi_q.wready), 
	.m_axi_bresp   (mem_reader_axi_q.bresp),  
	.m_axi_bvalid  (mem_reader_axi_q.bvalid), 
	.m_axi_bid     (mem_reader_axi_q.bid),
	.m_axi_bready  (mem_reader_axi_q.bready), 
	.m_axi_arid    (mem_reader_axi_q.arid), 
	.m_axi_araddr  (mem_reader_axi_q.araddr), 
	.m_axi_arlen   (mem_reader_axi_q.arlen), 
	.m_axi_arsize  (mem_reader_axi_q.arsize), 
	.m_axi_arvalid (mem_reader_axi_q.arvalid),
	.m_axi_arready (mem_reader_axi_q.arready),
	.m_axi_rid     (mem_reader_axi_q.rid),  
	.m_axi_rdata   (mem_reader_axi_q.rdata),  
	.m_axi_rresp   (mem_reader_axi_q.rresp),  
	.m_axi_rlast   (mem_reader_axi_q.rlast),  
	.m_axi_rvalid  (mem_reader_axi_q.rvalid), 
	.m_axi_rready  (mem_reader_axi_q.rready)
);



// AXI Crossbar: DMA_PCIS => DDR A/B/C/D
(* dont_touch = "true" *)
cl_axi_interconnect AXI_CROSSBAR
(
	.ACLK(clk),
	.ARESETN(slr_sync_aresetn),
	// DDR A
	.M00_AXI_araddr(ddr_a_pre.araddr),
	.M00_AXI_arburst(),
	.M00_AXI_arcache(),
	.M00_AXI_arid(ddr_a_pre.arid[6:0]),
	.M00_AXI_arlen(ddr_a_pre.arlen),
	.M00_AXI_arlock(),
	.M00_AXI_arprot(),
	.M00_AXI_arqos(),
	.M00_AXI_arready(ddr_a_pre.arready),
	.M00_AXI_arregion(),
	.M00_AXI_arsize(ddr_a_pre.arsize),
	.M00_AXI_arvalid(ddr_a_pre.arvalid),
	.M00_AXI_awaddr(ddr_a_pre.awaddr),
	.M00_AXI_awburst(),
	.M00_AXI_awcache(),
	.M00_AXI_awid(ddr_a_pre.awid[6:0]),
	.M00_AXI_awlen(ddr_a_pre.awlen),
	.M00_AXI_awlock(),
	.M00_AXI_awprot(),
	.M00_AXI_awqos(),
	.M00_AXI_awready(ddr_a_pre.awready),
	.M00_AXI_awregion(),
	.M00_AXI_awsize(ddr_a_pre.awsize),
	.M00_AXI_awvalid(ddr_a_pre.awvalid),
	.M00_AXI_bid(ddr_a_pre.bid[6:0]),
	.M00_AXI_bready(ddr_a_pre.bready),
	.M00_AXI_bresp(ddr_a_pre.bresp),
	.M00_AXI_bvalid(ddr_a_pre.bvalid),
	.M00_AXI_rdata(ddr_a_pre.rdata),
	.M00_AXI_rid(ddr_a_pre.rid[6:0]),
	.M00_AXI_rlast(ddr_a_pre.rlast),
	.M00_AXI_rready(ddr_a_pre.rready),
	.M00_AXI_rresp(ddr_a_pre.rresp),
	.M00_AXI_rvalid(ddr_a_pre.rvalid),
	.M00_AXI_wdata(ddr_a_pre.wdata),
	.M00_AXI_wlast(ddr_a_pre.wlast),
	.M00_AXI_wready(ddr_a_pre.wready),
	.M00_AXI_wstrb(ddr_a_pre.wstrb),
	.M00_AXI_wvalid(ddr_a_pre.wvalid),
	// DDR B
	.M01_AXI_araddr(ddr_b_pre.araddr),
	.M01_AXI_arburst(),
	.M01_AXI_arcache(),
	.M01_AXI_arid(ddr_b_pre.arid[6:0]),
	.M01_AXI_arlen(ddr_b_pre.arlen),
	.M01_AXI_arlock(),
	.M01_AXI_arprot(),
	.M01_AXI_arqos(),
	.M01_AXI_arready(ddr_b_pre.arready),
	.M01_AXI_arregion(),
	.M01_AXI_arsize(ddr_b_pre.arsize),
	.M01_AXI_arvalid(ddr_b_pre.arvalid),
	.M01_AXI_awaddr(ddr_b_pre.awaddr),
	.M01_AXI_awburst(),
	.M01_AXI_awcache(),
	.M01_AXI_awid(ddr_b_pre.awid[6:0]),
	.M01_AXI_awlen(ddr_b_pre.awlen),
	.M01_AXI_awlock(),
	.M01_AXI_awprot(),
	.M01_AXI_awqos(),
	.M01_AXI_awready(ddr_b_pre.awready),
	.M01_AXI_awregion(),
	.M01_AXI_awsize(ddr_b_pre.awsize),
	.M01_AXI_awvalid(ddr_b_pre.awvalid),
	.M01_AXI_bid(ddr_b_pre.bid[6:0]),
	.M01_AXI_bready(ddr_b_pre.bready),
	.M01_AXI_bresp(ddr_b_pre.bresp),
	.M01_AXI_bvalid(ddr_b_pre.bvalid),
	.M01_AXI_rdata(ddr_b_pre.rdata),
	.M01_AXI_rid(ddr_b_pre.rid[6:0]),
	.M01_AXI_rlast(ddr_b_pre.rlast),
	.M01_AXI_rready(ddr_b_pre.rready),
	.M01_AXI_rresp(ddr_b_pre.rresp),
	.M01_AXI_rvalid(ddr_b_pre.rvalid),
	.M01_AXI_wdata(ddr_b_pre.wdata),
	.M01_AXI_wlast(ddr_b_pre.wlast),
	.M01_AXI_wready(ddr_b_pre.wready),
	.M01_AXI_wstrb(ddr_b_pre.wstrb),
	.M01_AXI_wvalid(ddr_b_pre.wvalid),
	// DDR C
	.M02_AXI_araddr(ddr_c_pre.araddr),
	.M02_AXI_arburst(),
	.M02_AXI_arcache(),
	.M02_AXI_arid(ddr_c_pre.arid[6:0]),
	.M02_AXI_arlen(ddr_c_pre.arlen),
	.M02_AXI_arlock(),
	.M02_AXI_arprot(),
	.M02_AXI_arqos(),
	.M02_AXI_arready(ddr_c_pre.arready),
	.M02_AXI_arregion(),
	.M02_AXI_arsize(ddr_c_pre.arsize),
	.M02_AXI_arvalid(ddr_c_pre.arvalid),
	.M02_AXI_awaddr(ddr_c_pre.awaddr),
	.M02_AXI_awburst(),
	.M02_AXI_awcache(),
	.M02_AXI_awid(ddr_c_pre.awid[6:0]),
	.M02_AXI_awlen(ddr_c_pre.awlen),
	.M02_AXI_awlock(),
	.M02_AXI_awprot(),
	.M02_AXI_awqos(),
	.M02_AXI_awready(ddr_c_pre.awready),
	.M02_AXI_awregion(),
	.M02_AXI_awsize(ddr_c_pre.awsize),
	.M02_AXI_awvalid(ddr_c_pre.awvalid),
	.M02_AXI_bid(ddr_c_pre.bid[6:0]),
	.M02_AXI_bready(ddr_c_pre.bready),
	.M02_AXI_bresp(ddr_c_pre.bresp),
	.M02_AXI_bvalid(ddr_c_pre.bvalid),
	.M02_AXI_rdata(ddr_c_pre.rdata),
	.M02_AXI_rid(ddr_c_pre.rid[6:0]),
	.M02_AXI_rlast(ddr_c_pre.rlast),
	.M02_AXI_rready(ddr_c_pre.rready),
	.M02_AXI_rresp(ddr_c_pre.rresp),
	.M02_AXI_rvalid(ddr_c_pre.rvalid),
	.M02_AXI_wdata(ddr_c_pre.wdata),
	.M02_AXI_wlast(ddr_c_pre.wlast),
	.M02_AXI_wready(ddr_c_pre.wready),
	.M02_AXI_wstrb(ddr_c_pre.wstrb),
	.M02_AXI_wvalid(ddr_c_pre.wvalid),
	// DDR D
	.M03_AXI_araddr(ddr_d_pre.araddr),
	.M03_AXI_arburst(),
	.M03_AXI_arcache(),
	.M03_AXI_arid(ddr_d_pre.arid[6:0]),
	.M03_AXI_arlen(ddr_d_pre.arlen),
	.M03_AXI_arlock(),
	.M03_AXI_arprot(),
	.M03_AXI_arqos(),
	.M03_AXI_arready(ddr_d_pre.arready),
	.M03_AXI_arregion(),
	.M03_AXI_arsize(ddr_d_pre.arsize),
	.M03_AXI_arvalid(ddr_d_pre.arvalid),
	.M03_AXI_awaddr(ddr_d_pre.awaddr),
	.M03_AXI_awburst(),
	.M03_AXI_awcache(),
	.M03_AXI_awid(ddr_d_pre.awid[6:0]),
	.M03_AXI_awlen(ddr_d_pre.awlen),
	.M03_AXI_awlock(),
	.M03_AXI_awprot(),
	.M03_AXI_awqos(),
	.M03_AXI_awready(ddr_d_pre.awready),
	.M03_AXI_awregion(),
	.M03_AXI_awsize(ddr_d_pre.awsize),
	.M03_AXI_awvalid(ddr_d_pre.awvalid),
	.M03_AXI_bid(ddr_d_pre.bid[6:0]),
	.M03_AXI_bready(ddr_d_pre.bready),
	.M03_AXI_bresp(ddr_d_pre.bresp),
	.M03_AXI_bvalid(ddr_d_pre.bvalid),
	.M03_AXI_rdata(ddr_d_pre.rdata),
	.M03_AXI_rid(ddr_d_pre.rid[6:0]),
	.M03_AXI_rlast(ddr_d_pre.rlast),
	.M03_AXI_rready(ddr_d_pre.rready),
	.M03_AXI_rresp(ddr_d_pre.rresp),
	.M03_AXI_rvalid(ddr_d_pre.rvalid),
	.M03_AXI_wdata(ddr_d_pre.wdata),
	.M03_AXI_wlast(ddr_d_pre.wlast),
	.M03_AXI_wready(ddr_d_pre.wready),
	.M03_AXI_wstrb(ddr_d_pre.wstrb),
	.M03_AXI_wvalid(ddr_d_pre.wvalid),
	// DMA PCIS bus
	.S00_AXI_araddr({dma_pcis_bus_q.araddr[63:37], 1'b0, dma_pcis_bus_q.araddr[35:0]}),
	.S00_AXI_arburst(2'b1),
	.S00_AXI_arcache(4'b11),
	.S00_AXI_arid(dma_pcis_bus_q.arid[5:0]),
	.S00_AXI_arlen(dma_pcis_bus_q.arlen),
	.S00_AXI_arlock(1'b0),
	.S00_AXI_arprot(3'b10),
	.S00_AXI_arqos(4'b0),
	.S00_AXI_arready(dma_pcis_bus_q.arready),
	.S00_AXI_arregion(4'b0),
	.S00_AXI_arsize(dma_pcis_bus_q.arsize),
	.S00_AXI_arvalid(dma_pcis_bus_q.arvalid),
	.S00_AXI_awaddr({dma_pcis_bus_q.awaddr[63:37], 1'b0, dma_pcis_bus_q.awaddr[35:0]}),
	.S00_AXI_awburst(2'b1),
	.S00_AXI_awcache(4'b11),
	.S00_AXI_awid(dma_pcis_bus_q.awid[5:0]),
	.S00_AXI_awlen(dma_pcis_bus_q.awlen),
	.S00_AXI_awlock(1'b0),
	.S00_AXI_awprot(3'b10),
	.S00_AXI_awqos(4'b0),
	.S00_AXI_awready(dma_pcis_bus_q.awready),
	.S00_AXI_awregion(4'b0),
	.S00_AXI_awsize(dma_pcis_bus_q.awsize),
	.S00_AXI_awvalid(dma_pcis_bus_q.awvalid),
	.S00_AXI_bid(dma_pcis_bus_q.bid[5:0]),
	.S00_AXI_bready(dma_pcis_bus_q.bready),
	.S00_AXI_bresp(dma_pcis_bus_q.bresp),
	.S00_AXI_bvalid(dma_pcis_bus_q.bvalid),
	.S00_AXI_rdata(dma_pcis_bus_q.rdata),
	.S00_AXI_rid(dma_pcis_bus_q.rid[5:0]),
	.S00_AXI_rlast(dma_pcis_bus_q.rlast),
	.S00_AXI_rready(dma_pcis_bus_q.rready),
	.S00_AXI_rresp(dma_pcis_bus_q.rresp),
	.S00_AXI_rvalid(dma_pcis_bus_q.rvalid),
	.S00_AXI_wdata(dma_pcis_bus_q.wdata),
	.S00_AXI_wlast(dma_pcis_bus_q.wlast),
	.S00_AXI_wready(dma_pcis_bus_q.wready),
	.S00_AXI_wstrb(dma_pcis_bus_q.wstrb),
	.S00_AXI_wvalid(dma_pcis_bus_q.wvalid),
	// mem reader
	.S01_AXI_araddr({mem_reader_axi_q.araddr[63:37], 1'b0, mem_reader_axi_q.araddr[35:0]}),
	.S01_AXI_arburst(2'b1),
	.S01_AXI_arcache(4'b11),
	.S01_AXI_arid(mem_reader_axi_q.arid),
	.S01_AXI_arlen(mem_reader_axi_q.arlen),
	.S01_AXI_arlock(1'b0),
	.S01_AXI_arprot(3'b10),
	.S01_AXI_arqos(4'b0),
	.S01_AXI_arready(mem_reader_axi_q.arready),
	.S01_AXI_arregion(4'b0),
	.S01_AXI_arsize(mem_reader_axi_q.arsize),
	.S01_AXI_arvalid(mem_reader_axi_q.arvalid),
	.S01_AXI_awaddr({mem_reader_axi_q.awaddr[63:37], 1'b0, mem_reader_axi_q.awaddr[35:0]}),
	.S01_AXI_awburst(2'b1),
	.S01_AXI_awcache(4'b11),
	.S01_AXI_awid(mem_reader_axi_q.awid),
	.S01_AXI_awlen(mem_reader_axi_q.awlen),
	.S01_AXI_awlock(1'b0),
	.S01_AXI_awprot(3'b10),
	.S01_AXI_awqos(4'b0),
	.S01_AXI_awready(mem_reader_axi_q.awready),
	.S01_AXI_awregion(4'b0),
	.S01_AXI_awsize(mem_reader_axi_q.awsize),
	.S01_AXI_awvalid(mem_reader_axi_q.awvalid),
	.S01_AXI_bid(mem_reader_axi_q.bid),
	.S01_AXI_bready(mem_reader_axi_q.bready),
	.S01_AXI_bresp(mem_reader_axi_q.bresp),
	.S01_AXI_bvalid(mem_reader_axi_q.bvalid),
	.S01_AXI_rdata(mem_reader_axi_q.rdata),
	.S01_AXI_rid(mem_reader_axi_q.rid),
	.S01_AXI_rlast(mem_reader_axi_q.rlast),
	.S01_AXI_rready(mem_reader_axi_q.rready),
	.S01_AXI_rresp(mem_reader_axi_q.rresp),
	.S01_AXI_rvalid(mem_reader_axi_q.rvalid),
	.S01_AXI_wdata(mem_reader_axi_q.wdata),
	.S01_AXI_wlast(mem_reader_axi_q.wlast),
	.S01_AXI_wready(mem_reader_axi_q.wready),
	.S01_AXI_wstrb(mem_reader_axi_q.wstrb),
	.S01_AXI_wvalid(mem_reader_axi_q.wvalid)
);


// DDR A src -> dest path
src_register_slice DDR_A_SRC_SLICE (
	.aclk           (clk),
	.aresetn        (slr_sync_aresetn),
	// s
	.s_axi_awid     (ddr_a_pre.awid),
	.s_axi_awaddr   ({ddr_a_pre.awaddr[63:36], 2'b0, ddr_a_pre.awaddr[33:0]}),
	.s_axi_awlen    (ddr_a_pre.awlen),
	.s_axi_awsize   (ddr_a_pre.awsize),
	.s_axi_awburst  (2'b1),
	.s_axi_awlock   (1'b0),
	.s_axi_awcache  (4'b11),
	.s_axi_awprot   (3'b10),
	.s_axi_awregion (4'b0),
	.s_axi_awqos    (4'b0),
	.s_axi_awvalid  (ddr_a_pre.awvalid),
	.s_axi_awready  (ddr_a_pre.awready),
	.s_axi_wdata    (ddr_a_pre.wdata),
	.s_axi_wstrb    (ddr_a_pre.wstrb),
	.s_axi_wlast    (ddr_a_pre.wlast),
	.s_axi_wvalid   (ddr_a_pre.wvalid),
	.s_axi_wready   (ddr_a_pre.wready),
	.s_axi_bid      (ddr_a_pre.bid),
	.s_axi_bresp    (ddr_a_pre.bresp),
	.s_axi_bvalid   (ddr_a_pre.bvalid),
	.s_axi_bready   (ddr_a_pre.bready),
	.s_axi_arid     (ddr_a_pre.arid),
	.s_axi_araddr   ({ddr_a_pre.araddr[63:36], 2'b0, ddr_a_pre.araddr[33:0]}),
	.s_axi_arlen    (ddr_a_pre.arlen),
	.s_axi_arsize   (ddr_a_pre.arsize),
	.s_axi_arburst  (2'b1),
	.s_axi_arlock   (1'b0),
	.s_axi_arcache  (4'b11),
	.s_axi_arprot   (3'b10),
	.s_axi_arregion (4'b0),
	.s_axi_arqos    (4'b0),
	.s_axi_arvalid  (ddr_a_pre.arvalid),
	.s_axi_arready  (ddr_a_pre.arready),
	.s_axi_rid      (ddr_a_pre.rid),
	.s_axi_rdata    (ddr_a_pre.rdata),
	.s_axi_rresp    (ddr_a_pre.rresp),
	.s_axi_rlast    (ddr_a_pre.rlast),
	.s_axi_rvalid   (ddr_a_pre.rvalid),
	.s_axi_rready   (ddr_a_pre.rready),
	// m  
	.m_axi_awid     (ddr_a_src.awid),   
	.m_axi_awaddr   (ddr_a_src.awaddr), 
	.m_axi_awlen    (ddr_a_src.awlen),
	.m_axi_awsize   (ddr_a_src.awsize),
	.m_axi_awburst  (),
	.m_axi_awlock   (),
	.m_axi_awcache  (),
	.m_axi_awprot   (),
	.m_axi_awregion (),
	.m_axi_awqos    (),  
	.m_axi_awvalid  (ddr_a_src.awvalid),
	.m_axi_awready  (ddr_a_src.awready),
	.m_axi_wdata    (ddr_a_src.wdata),  
	.m_axi_wstrb    (ddr_a_src.wstrb),  
	.m_axi_wlast    (ddr_a_src.wlast),  
	.m_axi_wvalid   (ddr_a_src.wvalid), 
	.m_axi_wready   (ddr_a_src.wready), 
	.m_axi_bid      (ddr_a_src.bid),    
	.m_axi_bresp    (ddr_a_src.bresp),  
	.m_axi_bvalid   (ddr_a_src.bvalid), 
	.m_axi_bready   (ddr_a_src.bready), 
	.m_axi_arid     (ddr_a_src.arid),   
	.m_axi_araddr   (ddr_a_src.araddr), 
	.m_axi_arlen    (ddr_a_src.arlen),  
	.m_axi_arsize   (ddr_a_src.arsize),
	.m_axi_arburst  (),
	.m_axi_arlock   (),
	.m_axi_arcache  (),
	.m_axi_arprot   (),
	.m_axi_arregion (),
	.m_axi_arqos    (), 
	.m_axi_arvalid  (ddr_a_src.arvalid),
	.m_axi_arready  (ddr_a_src.arready),
	.m_axi_rid      (ddr_a_src.rid),    
	.m_axi_rdata    (ddr_a_src.rdata),  
	.m_axi_rresp    (ddr_a_src.rresp),  
	.m_axi_rlast    (ddr_a_src.rlast),  
	.m_axi_rvalid   (ddr_a_src.rvalid), 
	.m_axi_rready   (ddr_a_src.rready)
);

dest_register_slice DDR_A_DEST_SLICE
(
	.aclk           (clk),
	.aresetn        (slr_sync_aresetn),
	// s
	.s_axi_awid     (ddr_a_src.awid),
	.s_axi_awaddr   (ddr_a_src.awaddr),
	.s_axi_awlen    (ddr_a_src.awlen),
	.s_axi_awsize   (ddr_a_src.awsize),
	.s_axi_awburst  (2'b1),
	.s_axi_awlock   (1'b0),
	.s_axi_awcache  (4'b11),
	.s_axi_awprot   (3'b10),
	.s_axi_awregion (4'b0),
	.s_axi_awqos    (4'b0),
	.s_axi_awvalid  (ddr_a_src.awvalid),
	.s_axi_awready  (ddr_a_src.awready),
	.s_axi_wdata    (ddr_a_src.wdata),
	.s_axi_wstrb    (ddr_a_src.wstrb),
	.s_axi_wlast    (ddr_a_src.wlast),
	.s_axi_wvalid   (ddr_a_src.wvalid),
	.s_axi_wready   (ddr_a_src.wready),
	.s_axi_bid      (ddr_a_src.bid),
	.s_axi_bresp    (ddr_a_src.bresp),
	.s_axi_bvalid   (ddr_a_src.bvalid),
	.s_axi_bready   (ddr_a_src.bready),
	.s_axi_arid     (ddr_a_src.arid),
	.s_axi_araddr   (ddr_a_src.araddr),
	.s_axi_arlen    (ddr_a_src.arlen),
	.s_axi_arsize   (ddr_a_src.arsize),
	.s_axi_arburst  (2'b1),
	.s_axi_arlock   (1'b0),
	.s_axi_arcache  (4'b11),
	.s_axi_arprot   (3'b10),
	.s_axi_arregion (4'b0),
	.s_axi_arqos    (4'b0),
	.s_axi_arvalid  (ddr_a_src.arvalid),
	.s_axi_arready  (ddr_a_src.arready),
	.s_axi_rid      (ddr_a_src.rid),
	.s_axi_rdata    (ddr_a_src.rdata),
	.s_axi_rresp    (ddr_a_src.rresp),
	.s_axi_rlast    (ddr_a_src.rlast),
	.s_axi_rvalid   (ddr_a_src.rvalid),
	.s_axi_rready   (ddr_a_src.rready),
	// m
	.m_axi_awid     (ddr_a_dest.awid),   
	.m_axi_awaddr   (ddr_a_dest.awaddr), 
	.m_axi_awlen    (ddr_a_dest.awlen),
	.m_axi_awsize   (ddr_a_dest.awsize),
	.m_axi_awburst  (),
	.m_axi_awlock   (),
	.m_axi_awcache  (),
	.m_axi_awprot   (),
	.m_axi_awregion (),
	.m_axi_awqos    (),   
	.m_axi_awvalid  (ddr_a_dest.awvalid),
	.m_axi_awready  (ddr_a_dest.awready),
	.m_axi_wdata    (ddr_a_dest.wdata),  
	.m_axi_wstrb    (ddr_a_dest.wstrb),  
	.m_axi_wlast    (ddr_a_dest.wlast),  
	.m_axi_wvalid   (ddr_a_dest.wvalid), 
	.m_axi_wready   (ddr_a_dest.wready), 
	.m_axi_bid      (ddr_a_dest.bid),    
	.m_axi_bresp    (ddr_a_dest.bresp),  
	.m_axi_bvalid   (ddr_a_dest.bvalid), 
	.m_axi_bready   (ddr_a_dest.bready), 
	.m_axi_arid     (ddr_a_dest.arid),   
	.m_axi_araddr   (ddr_a_dest.araddr), 
	.m_axi_arlen    (ddr_a_dest.arlen),
	.m_axi_arsize   (ddr_a_dest.arsize),
	.m_axi_arburst  (),
	.m_axi_arlock   (),
	.m_axi_arcache  (),
	.m_axi_arprot   (),
	.m_axi_arregion (),
	.m_axi_arqos    (),   
	.m_axi_arvalid  (ddr_a_dest.arvalid),
	.m_axi_arready  (ddr_a_dest.arready),
	.m_axi_rid      (ddr_a_dest.rid),    
	.m_axi_rdata    (ddr_a_dest.rdata),  
	.m_axi_rresp    (ddr_a_dest.rresp),  
	.m_axi_rlast    (ddr_a_dest.rlast),  
	.m_axi_rvalid   (ddr_a_dest.rvalid), 
	.m_axi_rready   (ddr_a_dest.rready)
);

assign ddr_a_out.awid = {9'b0, ddr_a_dest.awid[6:0]};
assign ddr_a_out.awaddr = ddr_a_dest.awaddr;
assign ddr_a_out.awlen = ddr_a_dest.awlen;
assign ddr_a_out.awsize = ddr_a_dest.awsize;
assign ddr_a_out.awvalid = ddr_a_dest.awvalid;
assign ddr_a_dest.awready = ddr_a_out.awready;

assign ddr_a_out.wdata = ddr_a_dest.wdata;
assign ddr_a_out.wstrb = ddr_a_dest.wstrb;
assign ddr_a_out.wlast = ddr_a_dest.wlast;
assign ddr_a_out.wvalid = ddr_a_dest.wvalid;
assign ddr_a_dest.wready = ddr_a_out.wready;
assign ddr_a_out.wid = 16'b0;

assign ddr_a_dest.bid = {9'b0, ddr_a_out.bid[6:0]};
assign ddr_a_dest.bresp = ddr_a_out.bresp;
assign ddr_a_dest.bvalid = ddr_a_out.bvalid;
assign ddr_a_out.bready = ddr_a_dest.bready;

assign ddr_a_out.arid = {9'b0, ddr_a_dest.arid[6:0]};
assign ddr_a_out.araddr = ddr_a_dest.araddr;
assign ddr_a_out.arlen = ddr_a_dest.arlen;
assign ddr_a_out.arsize = ddr_a_dest.arsize;
assign ddr_a_out.arvalid = ddr_a_dest.arvalid;
assign ddr_a_dest.arready = ddr_a_out.arready;

assign ddr_a_dest.rid = {9'b0, ddr_a_out.rid[6:0]};
assign ddr_a_dest.rdata = ddr_a_out.rdata;
assign ddr_a_dest.rresp = ddr_a_out.rresp;
assign ddr_a_dest.rlast = ddr_a_out.rlast;
assign ddr_a_dest.rvalid = ddr_a_out.rvalid;
assign ddr_a_out.rready = ddr_a_dest.rready;

// DDR B src -> dest path
src_register_slice DDR_B_SRC_SLICE (
	.aclk           (clk),
	.aresetn        (slr_sync_aresetn),
	// s
	.s_axi_awid     (ddr_b_pre.awid),
	.s_axi_awaddr   ({ddr_b_pre.awaddr[63:36], 2'b0, ddr_b_pre.awaddr[33:0]}),
	.s_axi_awlen    (ddr_b_pre.awlen),
	.s_axi_awsize   (ddr_b_pre.awsize),
	.s_axi_awburst  (2'b1),
	.s_axi_awlock   (1'b0),
	.s_axi_awcache  (4'b11),
	.s_axi_awprot   (3'b10),
	.s_axi_awregion (4'b0),
	.s_axi_awqos    (4'b0),
	.s_axi_awvalid  (ddr_b_pre.awvalid),
	.s_axi_awready  (ddr_b_pre.awready),
	.s_axi_wdata    (ddr_b_pre.wdata),
	.s_axi_wstrb    (ddr_b_pre.wstrb),
	.s_axi_wlast    (ddr_b_pre.wlast),
	.s_axi_wvalid   (ddr_b_pre.wvalid),
	.s_axi_wready   (ddr_b_pre.wready),
	.s_axi_bid      (ddr_b_pre.bid),
	.s_axi_bresp    (ddr_b_pre.bresp),
	.s_axi_bvalid   (ddr_b_pre.bvalid),
	.s_axi_bready   (ddr_b_pre.bready),
	.s_axi_arid     (ddr_b_pre.arid),
	.s_axi_araddr   ({ddr_b_pre.araddr[63:36], 2'b0, ddr_b_pre.araddr[33:0]}),
	.s_axi_arlen    (ddr_b_pre.arlen),
	.s_axi_arsize   (ddr_b_pre.arsize),
	.s_axi_arburst  (2'b1),
	.s_axi_arlock   (1'b0),
	.s_axi_arcache  (4'b11),
	.s_axi_arprot   (3'b10),
	.s_axi_arregion (4'b0),
	.s_axi_arqos    (4'b0),
	.s_axi_arvalid  (ddr_b_pre.arvalid),
	.s_axi_arready  (ddr_b_pre.arready),
	.s_axi_rid      (ddr_b_pre.rid),
	.s_axi_rdata    (ddr_b_pre.rdata),
	.s_axi_rresp    (ddr_b_pre.rresp),
	.s_axi_rlast    (ddr_b_pre.rlast),
	.s_axi_rvalid   (ddr_b_pre.rvalid),
	.s_axi_rready   (ddr_b_pre.rready),
	// m  
	.m_axi_awid     (ddr_b_src.awid),   
	.m_axi_awaddr   (ddr_b_src.awaddr), 
	.m_axi_awlen    (ddr_b_src.awlen),
	.m_axi_awsize   (ddr_b_src.awsize),
	.m_axi_awburst  (),
	.m_axi_awlock   (),
	.m_axi_awcache  (),
	.m_axi_awprot   (),
	.m_axi_awregion (),
	.m_axi_awqos    (),  
	.m_axi_awvalid  (ddr_b_src.awvalid),
	.m_axi_awready  (ddr_b_src.awready),
	.m_axi_wdata    (ddr_b_src.wdata),  
	.m_axi_wstrb    (ddr_b_src.wstrb),  
	.m_axi_wlast    (ddr_b_src.wlast),  
	.m_axi_wvalid   (ddr_b_src.wvalid), 
	.m_axi_wready   (ddr_b_src.wready), 
	.m_axi_bid      (ddr_b_src.bid),    
	.m_axi_bresp    (ddr_b_src.bresp),  
	.m_axi_bvalid   (ddr_b_src.bvalid), 
	.m_axi_bready   (ddr_b_src.bready), 
	.m_axi_arid     (ddr_b_src.arid),   
	.m_axi_araddr   (ddr_b_src.araddr), 
	.m_axi_arlen    (ddr_b_src.arlen),  
	.m_axi_arsize   (ddr_b_src.arsize),
	.m_axi_arburst  (),
	.m_axi_arlock   (),
	.m_axi_arcache  (),
	.m_axi_arprot   (),
	.m_axi_arregion (),
	.m_axi_arqos    (), 
	.m_axi_arvalid  (ddr_b_src.arvalid),
	.m_axi_arready  (ddr_b_src.arready),
	.m_axi_rid      (ddr_b_src.rid),    
	.m_axi_rdata    (ddr_b_src.rdata),  
	.m_axi_rresp    (ddr_b_src.rresp),  
	.m_axi_rlast    (ddr_b_src.rlast),  
	.m_axi_rvalid   (ddr_b_src.rvalid), 
	.m_axi_rready   (ddr_b_src.rready)
);

dest_register_slice DDR_B_DEST_SLICE
(
	.aclk           (clk),
	.aresetn        (slr_sync_aresetn),
	// s
	.s_axi_awid     (ddr_b_src.awid),
	.s_axi_awaddr   (ddr_b_src.awaddr),
	.s_axi_awlen    (ddr_b_src.awlen),
	.s_axi_awsize   (ddr_b_src.awsize),
	.s_axi_awburst  (2'b1),
	.s_axi_awlock   (1'b0),
	.s_axi_awcache  (4'b11),
	.s_axi_awprot   (3'b10),
	.s_axi_awregion (4'b0),
	.s_axi_awqos    (4'b0),
	.s_axi_awvalid  (ddr_b_src.awvalid),
	.s_axi_awready  (ddr_b_src.awready),
	.s_axi_wdata    (ddr_b_src.wdata),
	.s_axi_wstrb    (ddr_b_src.wstrb),
	.s_axi_wlast    (ddr_b_src.wlast),
	.s_axi_wvalid   (ddr_b_src.wvalid),
	.s_axi_wready   (ddr_b_src.wready),
	.s_axi_bid      (ddr_b_src.bid),
	.s_axi_bresp    (ddr_b_src.bresp),
	.s_axi_bvalid   (ddr_b_src.bvalid),
	.s_axi_bready   (ddr_b_src.bready),
	.s_axi_arid     (ddr_b_src.arid),
	.s_axi_araddr   (ddr_b_src.araddr),
	.s_axi_arlen    (ddr_b_src.arlen),
	.s_axi_arsize   (ddr_b_src.arsize),
	.s_axi_arburst  (2'b1),
	.s_axi_arlock   (1'b0),
	.s_axi_arcache  (4'b11),
	.s_axi_arprot   (3'b10),
	.s_axi_arregion (4'b0),
	.s_axi_arqos    (4'b0),
	.s_axi_arvalid  (ddr_b_src.arvalid),
	.s_axi_arready  (ddr_b_src.arready),
	.s_axi_rid      (ddr_b_src.rid),
	.s_axi_rdata    (ddr_b_src.rdata),
	.s_axi_rresp    (ddr_b_src.rresp),
	.s_axi_rlast    (ddr_b_src.rlast),
	.s_axi_rvalid   (ddr_b_src.rvalid),
	.s_axi_rready   (ddr_b_src.rready),
	// m
	.m_axi_awid     (ddr_b_dest.awid),   
	.m_axi_awaddr   (ddr_b_dest.awaddr), 
	.m_axi_awlen    (ddr_b_dest.awlen),
	.m_axi_awsize   (ddr_b_dest.awsize),
	.m_axi_awburst  (),
	.m_axi_awlock   (),
	.m_axi_awcache  (),
	.m_axi_awprot   (),
	.m_axi_awregion (),
	.m_axi_awqos    (),   
	.m_axi_awvalid  (ddr_b_dest.awvalid),
	.m_axi_awready  (ddr_b_dest.awready),
	.m_axi_wdata    (ddr_b_dest.wdata),  
	.m_axi_wstrb    (ddr_b_dest.wstrb),  
	.m_axi_wlast    (ddr_b_dest.wlast),  
	.m_axi_wvalid   (ddr_b_dest.wvalid), 
	.m_axi_wready   (ddr_b_dest.wready), 
	.m_axi_bid      (ddr_b_dest.bid),    
	.m_axi_bresp    (ddr_b_dest.bresp),  
	.m_axi_bvalid   (ddr_b_dest.bvalid), 
	.m_axi_bready   (ddr_b_dest.bready), 
	.m_axi_arid     (ddr_b_dest.arid),   
	.m_axi_araddr   (ddr_b_dest.araddr), 
	.m_axi_arlen    (ddr_b_dest.arlen),
	.m_axi_arsize   (ddr_b_dest.arsize),
	.m_axi_arburst  (),
	.m_axi_arlock   (),
	.m_axi_arcache  (),
	.m_axi_arprot   (),
	.m_axi_arregion (),
	.m_axi_arqos    (),   
	.m_axi_arvalid  (ddr_b_dest.arvalid),
	.m_axi_arready  (ddr_b_dest.arready),
	.m_axi_rid      (ddr_b_dest.rid),    
	.m_axi_rdata    (ddr_b_dest.rdata),  
	.m_axi_rresp    (ddr_b_dest.rresp),  
	.m_axi_rlast    (ddr_b_dest.rlast),  
	.m_axi_rvalid   (ddr_b_dest.rvalid), 
	.m_axi_rready   (ddr_b_dest.rready)
);

assign ddr_b_out.awid = {9'b0, ddr_b_dest.awid[6:0]};
assign ddr_b_out.awaddr = ddr_b_dest.awaddr;
assign ddr_b_out.awlen = ddr_b_dest.awlen;
assign ddr_b_out.awsize = ddr_b_dest.awsize;
assign ddr_b_out.awvalid = ddr_b_dest.awvalid;
assign ddr_b_dest.awready = ddr_b_out.awready;

assign ddr_b_out.wdata = ddr_b_dest.wdata;
assign ddr_b_out.wstrb = ddr_b_dest.wstrb;
assign ddr_b_out.wlast = ddr_b_dest.wlast;
assign ddr_b_out.wvalid = ddr_b_dest.wvalid;
assign ddr_b_dest.wready = ddr_b_out.wready;
assign ddr_b_out.wid = 16'b0;

assign ddr_b_dest.bid = {9'b0, ddr_b_out.bid[6:0]};
assign ddr_b_dest.bresp = ddr_b_out.bresp;
assign ddr_b_dest.bvalid = ddr_b_out.bvalid;
assign ddr_b_out.bready = ddr_b_dest.bready;

assign ddr_b_out.arid = {9'b0, ddr_b_dest.arid[6:0]};
assign ddr_b_out.araddr = ddr_b_dest.araddr;
assign ddr_b_out.arlen = ddr_b_dest.arlen;
assign ddr_b_out.arsize = ddr_b_dest.arsize;
assign ddr_b_out.arvalid = ddr_b_dest.arvalid;
assign ddr_b_dest.arready = ddr_b_out.arready;

assign ddr_b_dest.rid = {9'b0, ddr_b_out.rid[6:0]};
assign ddr_b_dest.rdata = ddr_b_out.rdata;
assign ddr_b_dest.rresp = ddr_b_out.rresp;
assign ddr_b_dest.rlast = ddr_b_out.rlast;
assign ddr_b_dest.rvalid = ddr_b_out.rvalid;
assign ddr_b_out.rready = ddr_b_dest.rready;


// DDR D src -> dest path
src_register_slice DDR_D_SRC_SLICE (
	.aclk           (clk),
	.aresetn        (slr_sync_aresetn),
	// s
	.s_axi_awid     (ddr_d_pre.awid),
	.s_axi_awaddr   ({ddr_d_pre.awaddr[63:36], 2'b0, ddr_d_pre.awaddr[33:0]}),
	.s_axi_awlen    (ddr_d_pre.awlen),
	.s_axi_awsize   (ddr_d_pre.awsize),
	.s_axi_awburst  (2'b1),
	.s_axi_awlock   (1'b0),
	.s_axi_awcache  (4'b11),
	.s_axi_awprot   (3'b10),
	.s_axi_awregion (4'b0),
	.s_axi_awqos    (4'b0),
	.s_axi_awvalid  (ddr_d_pre.awvalid),
	.s_axi_awready  (ddr_d_pre.awready),
	.s_axi_wdata    (ddr_d_pre.wdata),
	.s_axi_wstrb    (ddr_d_pre.wstrb),
	.s_axi_wlast    (ddr_d_pre.wlast),
	.s_axi_wvalid   (ddr_d_pre.wvalid),
	.s_axi_wready   (ddr_d_pre.wready),
	.s_axi_bid      (ddr_d_pre.bid),
	.s_axi_bresp    (ddr_d_pre.bresp),
	.s_axi_bvalid   (ddr_d_pre.bvalid),
	.s_axi_bready   (ddr_d_pre.bready),
	.s_axi_arid     (ddr_d_pre.arid),
	.s_axi_araddr   ({ddr_d_pre.araddr[63:36], 2'b0, ddr_d_pre.araddr[33:0]}),
	.s_axi_arlen    (ddr_d_pre.arlen),
	.s_axi_arsize   (ddr_d_pre.arsize),
	.s_axi_arburst  (2'b1),
	.s_axi_arlock   (1'b0),
	.s_axi_arcache  (4'b11),
	.s_axi_arprot   (3'b10),
	.s_axi_arregion (4'b0),
	.s_axi_arqos    (4'b0),
	.s_axi_arvalid  (ddr_d_pre.arvalid),
	.s_axi_arready  (ddr_d_pre.arready),
	.s_axi_rid      (ddr_d_pre.rid),
	.s_axi_rdata    (ddr_d_pre.rdata),
	.s_axi_rresp    (ddr_d_pre.rresp),
	.s_axi_rlast    (ddr_d_pre.rlast),
	.s_axi_rvalid   (ddr_d_pre.rvalid),
	.s_axi_rready   (ddr_d_pre.rready),
	// m  
	.m_axi_awid     (ddr_d_src.awid),   
	.m_axi_awaddr   (ddr_d_src.awaddr), 
	.m_axi_awlen    (ddr_d_src.awlen),
	.m_axi_awsize   (ddr_d_src.awsize),
	.m_axi_awburst  (),
	.m_axi_awlock   (),
	.m_axi_awcache  (),
	.m_axi_awprot   (),
	.m_axi_awregion (),
	.m_axi_awqos    (),  
	.m_axi_awvalid  (ddr_d_src.awvalid),
	.m_axi_awready  (ddr_d_src.awready),
	.m_axi_wdata    (ddr_d_src.wdata),  
	.m_axi_wstrb    (ddr_d_src.wstrb),  
	.m_axi_wlast    (ddr_d_src.wlast),  
	.m_axi_wvalid   (ddr_d_src.wvalid), 
	.m_axi_wready   (ddr_d_src.wready), 
	.m_axi_bid      (ddr_d_src.bid),    
	.m_axi_bresp    (ddr_d_src.bresp),  
	.m_axi_bvalid   (ddr_d_src.bvalid), 
	.m_axi_bready   (ddr_d_src.bready), 
	.m_axi_arid     (ddr_d_src.arid),   
	.m_axi_araddr   (ddr_d_src.araddr), 
	.m_axi_arlen    (ddr_d_src.arlen),  
	.m_axi_arsize   (ddr_d_src.arsize),
	.m_axi_arburst  (),
	.m_axi_arlock   (),
	.m_axi_arcache  (),
	.m_axi_arprot   (),
	.m_axi_arregion (),
	.m_axi_arqos    (), 
	.m_axi_arvalid  (ddr_d_src.arvalid),
	.m_axi_arready  (ddr_d_src.arready),
	.m_axi_rid      (ddr_d_src.rid),    
	.m_axi_rdata    (ddr_d_src.rdata),  
	.m_axi_rresp    (ddr_d_src.rresp),  
	.m_axi_rlast    (ddr_d_src.rlast),  
	.m_axi_rvalid   (ddr_d_src.rvalid), 
	.m_axi_rready   (ddr_d_src.rready)
);

dest_register_slice DDR_D_DEST_SLICE
(
	.aclk           (clk),
	.aresetn        (slr_sync_aresetn),
	// s
	.s_axi_awid     (ddr_d_src.awid),
	.s_axi_awaddr   (ddr_d_src.awaddr),
	.s_axi_awlen    (ddr_d_src.awlen),
	.s_axi_awsize   (ddr_d_src.awsize),
	.s_axi_awburst  (2'b1),
	.s_axi_awlock   (1'b0),
	.s_axi_awcache  (4'b11),
	.s_axi_awprot   (3'b10),
	.s_axi_awregion (4'b0),
	.s_axi_awqos    (4'b0),
	.s_axi_awvalid  (ddr_d_src.awvalid),
	.s_axi_awready  (ddr_d_src.awready),
	.s_axi_wdata    (ddr_d_src.wdata),
	.s_axi_wstrb    (ddr_d_src.wstrb),
	.s_axi_wlast    (ddr_d_src.wlast),
	.s_axi_wvalid   (ddr_d_src.wvalid),
	.s_axi_wready   (ddr_d_src.wready),
	.s_axi_bid      (ddr_d_src.bid),
	.s_axi_bresp    (ddr_d_src.bresp),
	.s_axi_bvalid   (ddr_d_src.bvalid),
	.s_axi_bready   (ddr_d_src.bready),
	.s_axi_arid     (ddr_d_src.arid),
	.s_axi_araddr   (ddr_d_src.araddr),
	.s_axi_arlen    (ddr_d_src.arlen),
	.s_axi_arsize   (ddr_d_src.arsize),
	.s_axi_arburst  (2'b1),
	.s_axi_arlock   (1'b0),
	.s_axi_arcache  (4'b11),
	.s_axi_arprot   (3'b10),
	.s_axi_arregion (4'b0),
	.s_axi_arqos    (4'b0),
	.s_axi_arvalid  (ddr_d_src.arvalid),
	.s_axi_arready  (ddr_d_src.arready),
	.s_axi_rid      (ddr_d_src.rid),
	.s_axi_rdata    (ddr_d_src.rdata),
	.s_axi_rresp    (ddr_d_src.rresp),
	.s_axi_rlast    (ddr_d_src.rlast),
	.s_axi_rvalid   (ddr_d_src.rvalid),
	.s_axi_rready   (ddr_d_src.rready),
	// m
	.m_axi_awid     (ddr_d_dest.awid),   
	.m_axi_awaddr   (ddr_d_dest.awaddr), 
	.m_axi_awlen    (ddr_d_dest.awlen),
	.m_axi_awsize   (ddr_d_dest.awsize),
	.m_axi_awburst  (),
	.m_axi_awlock   (),
	.m_axi_awcache  (),
	.m_axi_awprot   (),
	.m_axi_awregion (),
	.m_axi_awqos    (),   
	.m_axi_awvalid  (ddr_d_dest.awvalid),
	.m_axi_awready  (ddr_d_dest.awready),
	.m_axi_wdata    (ddr_d_dest.wdata),  
	.m_axi_wstrb    (ddr_d_dest.wstrb),  
	.m_axi_wlast    (ddr_d_dest.wlast),  
	.m_axi_wvalid   (ddr_d_dest.wvalid), 
	.m_axi_wready   (ddr_d_dest.wready), 
	.m_axi_bid      (ddr_d_dest.bid),    
	.m_axi_bresp    (ddr_d_dest.bresp),  
	.m_axi_bvalid   (ddr_d_dest.bvalid), 
	.m_axi_bready   (ddr_d_dest.bready), 
	.m_axi_arid     (ddr_d_dest.arid),   
	.m_axi_araddr   (ddr_d_dest.araddr), 
	.m_axi_arlen    (ddr_d_dest.arlen),
	.m_axi_arsize   (ddr_d_dest.arsize),
	.m_axi_arburst  (),
	.m_axi_arlock   (),
	.m_axi_arcache  (),
	.m_axi_arprot   (),
	.m_axi_arregion (),
	.m_axi_arqos    (),   
	.m_axi_arvalid  (ddr_d_dest.arvalid),
	.m_axi_arready  (ddr_d_dest.arready),
	.m_axi_rid      (ddr_d_dest.rid),    
	.m_axi_rdata    (ddr_d_dest.rdata),  
	.m_axi_rresp    (ddr_d_dest.rresp),  
	.m_axi_rlast    (ddr_d_dest.rlast),  
	.m_axi_rvalid   (ddr_d_dest.rvalid), 
	.m_axi_rready   (ddr_d_dest.rready)
);

assign ddr_d_out.awid = {9'b0, ddr_d_dest.awid[6:0]};
assign ddr_d_out.awaddr = ddr_d_dest.awaddr;
assign ddr_d_out.awlen = ddr_d_dest.awlen;
assign ddr_d_out.awsize = ddr_d_dest.awsize;
assign ddr_d_out.awvalid = ddr_d_dest.awvalid;
assign ddr_d_dest.awready = ddr_d_out.awready;

assign ddr_d_out.wdata = ddr_d_dest.wdata;
assign ddr_d_out.wstrb = ddr_d_dest.wstrb;
assign ddr_d_out.wlast = ddr_d_dest.wlast;
assign ddr_d_out.wvalid = ddr_d_dest.wvalid;
assign ddr_d_dest.wready = ddr_d_out.wready;
assign ddr_d_out.wid = 16'b0;

assign ddr_d_dest.bid = {9'b0, ddr_d_out.bid[6:0]};
assign ddr_d_dest.bresp = ddr_d_out.bresp;
assign ddr_d_dest.bvalid = ddr_d_out.bvalid;
assign ddr_d_out.bready = ddr_d_dest.bready;

assign ddr_d_out.arid = {9'b0, ddr_d_dest.arid[6:0]};
assign ddr_d_out.araddr = ddr_d_dest.araddr;
assign ddr_d_out.arlen = ddr_d_dest.arlen;
assign ddr_d_out.arsize = ddr_d_dest.arsize;
assign ddr_d_out.arvalid = ddr_d_dest.arvalid;
assign ddr_d_dest.arready = ddr_d_out.arready;

assign ddr_d_dest.rid = {9'b0, ddr_d_out.rid[6:0]};
assign ddr_d_dest.rdata = ddr_d_out.rdata;
assign ddr_d_dest.rresp = ddr_d_out.rresp;
assign ddr_d_dest.rlast = ddr_d_out.rlast;
assign ddr_d_dest.rvalid = ddr_d_out.rvalid;
assign ddr_d_out.rready = ddr_d_dest.rready;

// DDR C
axi_register_slice DDR_C_TST_AXI4_REG_SLC (
	.aclk           (clk),
	.aresetn        (slr_sync_aresetn),
	// s                                                                                               
	.s_axi_awid     (ddr_c_pre.awid),
	.s_axi_awaddr   ({ddr_c_pre.awaddr[63:36], 2'b0, ddr_c_pre.awaddr[33:0]}),
	.s_axi_awlen    (ddr_c_pre.awlen),
	.s_axi_awsize   (ddr_c_pre.awsize),
	.s_axi_awvalid  (ddr_c_pre.awvalid),
	.s_axi_awready  (ddr_c_pre.awready),
	.s_axi_wdata    (ddr_c_pre.wdata),
	.s_axi_wstrb    (ddr_c_pre.wstrb),
	.s_axi_wlast    (ddr_c_pre.wlast),
	.s_axi_wvalid   (ddr_c_pre.wvalid),
	.s_axi_wready   (ddr_c_pre.wready),
	.s_axi_bid      (ddr_c_pre.bid),
	.s_axi_bresp    (ddr_c_pre.bresp),
	.s_axi_bvalid   (ddr_c_pre.bvalid),
	.s_axi_bready   (ddr_c_pre.bready),
	.s_axi_arid     (ddr_c_pre.arid),
	.s_axi_araddr   ({ddr_c_pre.araddr[63:36], 2'b0, ddr_c_pre.araddr[33:0]}),
	.s_axi_arlen    (ddr_c_pre.arlen),
	.s_axi_arsize   (ddr_c_pre.arsize),
	.s_axi_arvalid  (ddr_c_pre.arvalid),
	.s_axi_arready  (ddr_c_pre.arready),
	.s_axi_rid      (ddr_c_pre.rid),
	.s_axi_rdata    (ddr_c_pre.rdata),
	.s_axi_rresp    (ddr_c_pre.rresp),
	.s_axi_rlast    (ddr_c_pre.rlast),
	.s_axi_rvalid   (ddr_c_pre.rvalid),
	.s_axi_rready   (ddr_c_pre.rready),
	// m
	.m_axi_awid     (ddr_c_out.awid),   
	.m_axi_awaddr   (ddr_c_out.awaddr), 
	.m_axi_awlen    (ddr_c_out.awlen),  
	.m_axi_awsize   (ddr_c_out.awsize),
	.m_axi_awvalid  (ddr_c_out.awvalid),
	.m_axi_awready  (ddr_c_out.awready),
	.m_axi_wdata    (ddr_c_out.wdata),  
	.m_axi_wstrb    (ddr_c_out.wstrb),  
	.m_axi_wlast    (ddr_c_out.wlast),  
	.m_axi_wvalid   (ddr_c_out.wvalid), 
	.m_axi_wready   (ddr_c_out.wready), 
	.m_axi_bid      (ddr_c_out.bid),    
	.m_axi_bresp    (ddr_c_out.bresp),  
	.m_axi_bvalid   (ddr_c_out.bvalid), 
	.m_axi_bready   (ddr_c_out.bready), 
	.m_axi_arid     (ddr_c_out.arid),   
	.m_axi_araddr   (ddr_c_out.araddr), 
	.m_axi_arlen    (ddr_c_out.arlen),  
	.m_axi_arsize   (ddr_c_out.arsize),
	.m_axi_arvalid  (ddr_c_out.arvalid),
	.m_axi_arready  (ddr_c_out.arready),
	.m_axi_rid      (ddr_c_out.rid),    
	.m_axi_rdata    (ddr_c_out.rdata),  
	.m_axi_rresp    (ddr_c_out.rresp),  
	.m_axi_rlast    (ddr_c_out.rlast),  
	.m_axi_rvalid   (ddr_c_out.rvalid), 
	.m_axi_rready   (ddr_c_out.rready)
);



endmodule

