`ifndef CL_DRAM_PERF_DEFINES
`define CL_DRAM_PERF_DEFINES

`define CL_NAME cl_dram_perf
`define FPGA_LESS_RST

`endif
